`timescale 1ps/1ps

module OP#(
   parameter XLEN = 32  
)(
    input    [XLEN-1:0]  op_data_1,
    input    [XLEN-1:0]  op_data_2,
    output   [XLEN-1:0]  op_result
);
    



endmodule